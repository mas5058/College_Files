library verilog;
use verilog.vl_types.all;
entity hw7_1_vlg_vec_tst is
end hw7_1_vlg_vec_tst;
