-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--Michael Sarlo
--lab 1
--8/30/16
--xor gate
---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
entity xor2
        port(a, b : in std_logic
             z    : out std_logic)
    end xor2


architecture arch of xor2 is
begin
    z <= a xor b
end arch;