-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--Michael Sarlo
--lab 1
--8/23/16
--single bit adder
-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
library ieee
use ieee.std_logic_1164.all;
entity adder is
    port{
    a     : in std_logic_vector(32 downto 0);
    b       : in std_logic;
    c       : out std_logic;
    };

    
    
    1 
    2 
    3 
    4 
    5 
    6 
    7 
    8 
    9 
    10
    11