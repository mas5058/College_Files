library verilog;
use verilog.vl_types.all;
entity hw6_vlg_check_tst is
    port(
        q               : in     vl_logic;
        qn              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end hw6_vlg_check_tst;
