-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--Michael Sarlo
--lab 1
--8/30/16
--or gate
---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------

entity or3
        port(a, b, c : in std_logic
             z    : out std_logic)
    end or3


architecture arch of or3 is
begin
    z <= a or b or c;
end arch;