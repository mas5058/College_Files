library verilog;
use verilog.vl_types.all;
entity hw6_vlg_vec_tst is
end hw6_vlg_vec_tst;
