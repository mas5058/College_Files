entity receive
	port(input : in std_logic_vector(15 downto 0);
		  
		  )